//this module implements an N-bit ripple carry adder

